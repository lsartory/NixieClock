library ieee;
use ieee.std_logic_1164.all;

entity Nixie is
	port
	(
		CLK : in std_logic
	);
end Nixie;


architecture Nixie_Arch of Nixie is
begin

end architecture;
